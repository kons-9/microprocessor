`timescale 1ns / 1ps

`include "define.v"

module forwarding(
    input wire reg1_addrEW,
    input wire reg2_addrEW,
    input wire dst_reg_data;

    output wire reg1_data,
    output wire reg2_data,
    output wire reg1_signal,
    output wire reg2_sig
    );

    




endmodule